LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY REG IS
PORT(
	REG_CLK: IN STD_LOGIC;
	A_IN: IN STD_LOGIC;
	A_OUT: IN STD_LOGIC;
	INPUT_DATA: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	OUTPUT_DATA:  OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	OUTPUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	
);
END REG;


ARCHITECTURE REG OF REG IS 

BEGIN

PROCESS(REG_CLK,A_OUT)
VARIABLE DATA: STD_LOGIC_VECTOR(7 DOWNTO 0);
VARIABLE OUT_DATA: STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
IF(A_OUT='1') THEN
	OUT_DATA:=DATA;
ELSE IF(A_OUT='0') THEN
	OUT_DATA:="ZZZZZZZZ";
END IF;
END IF;

IF(REG_CLK'EVENT AND REG_CLK='1') THEN
	IF(A_IN='1') THEN
		DATA:= INPUT_DATA;
		

	END IF;
	
	OUTPUT_DATA<=OUT_DATA;
END IF;
IF(REG_CLK'EVENT AND REG_CLK='0') THEN
	IF(A_IN='1') THEN
		
		OUTPUT<=INPUT_DATA;

	END IF;
	
	
END IF;

END PROCESS;

END REG;

	

		
		