LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


ENTITY RAM IS
PORT(
	ADDRESS: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	DATA_IN: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	DATA_OUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	RAM_IN: IN STD_LOGIC;
	RAM_OUT: IN STD_LOGIC;
	RAM_CLK: IN STD_LOGIC;
	ADDRESS_IN:IN STD_LOGIC

);
END RAM;

ARCHITECTURE RAM OF RAM IS

TYPE MEMORY IS ARRAY (0 TO 15) OF STD_LOGIC_VECTOR(7 DOWNTO 0);

SIGNAL RANDOM_MEMORY: MEMORY:=(
					"00001001",--0
					"00011010",--1
					"00101101",--2
					"00000000",--3
					"00000000",--4
					"00000000",--5
					"00000000",--6
					"00000000",--7
					"00000000",--8
					"00000010",--9
					"00000010",--10
					"00000000",--11
					"00000000",--12
					"00000000",--13
					"00000000",--14
					"00000000" --15
				);
					
BEGIN

PROCESS(RAM_CLK,RAM_IN,RAM_OUT)
VARIABLE DATA: STD_LOGIC_VECTOR(7 DOWNTO 0);
VARIABLE ADDRESS_BUFFER:STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
IF(ADDRESS_IN='1') THEN
ADDRESS_BUFFER:=ADDRESS;
END IF;

IF (RAM_OUT='1') THEN
	DATA:=RANDOM_MEMORY(CONV_INTEGER(ADDRESS_BUFFER));
ELSE IF (RAM_OUT='0') THEN 
	DATA:="ZZZZZZZZ";
END IF;
END IF;

IF(RAM_CLK'EVENT AND RAM_CLK='0') THEN
	IF(RAM_IN='1') THEN
		RANDOM_MEMORY(CONV_INTEGER(ADDRESS_BUFFER))<=DATA_IN;
	END IF;
END IF;
IF(RAM_CLK'EVENT AND RAM_CLK='1') THEN
	
DATA_OUT<=DATA;


END IF;
END PROCESS;
END RAM;