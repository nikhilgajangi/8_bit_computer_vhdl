LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CONTROL_UNIT IS
PORT( 
	CONTROL_BITS: OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
	CU_CLK: IN STD_LOGIC;
	OPCODE: IN STD_LOGIC_VECTOR(3 DOWNTO 0)
);
END CONTROL_UNIT;

ARCHITECTURE CONTROL_UNIT OF CONTROL_UNIT IS
SIGNAL STEP: STD_LOGIC_VECTOR(2 DOWNTO 0):="000";
SIGNAL ADDRESS: STD_LOGIC_VECTOR(6 DOWNTO 0);
TYPE CONTROL_MEMORY IS ARRAY(0 TO 59) OF STD_LOGIC_VECTOR(12 DOWNTO 0);

                                    --    PC_OUT,PC_INC,ID_IN,ID_OUT,ARITH_SELECT,ALU_OUT,A_IN,A_OUT,B_IN,B_OUT,RAM_IN,RAM_OUT,ADD_IN),
					
CONSTANT CONTROL_DATA: CONTROL_MEMORY:= (
						"1000000000001",--0
						"0110000000010",--1
						"0001000000001",--2
						"0000001000010",--3
						"0000000000000",--4
						"0000000000000",--5
						"0000000000000",--6
						"0000000000000",--7
						"0000000000000",--8
						"0000000000000",--9
						"0001000000001",--10
						"0000000010010",--11
						"0000000000000",--12
						"0000000000000",--13
						"0000000000000",--14
						"0000000000000",--15
						"0000000000000",--16
						"0000000000000",--17
						"0001100000001",--18
						"0000010000100",--19
						"0000000000000",--20
						"0000000000000",--21
						"0000000000000",--22
						"0000000000000",--23
						"0000000000000",--24
						"0000000000000",--25
						"0001000000001",--26
						"0000010000100",--27
						"0000000000000",--28
						"0000000000000",--29
						"0000000000000",--30
						"0000000000000",--31
						"0000000000000",--32
						"0000000000000",--33
						"0000000000000",--34
						"0000000000000",--35
						"0000000000000",--36
						"0000000000000",--37
						"0000000000000",--38
						"0000000000000",--39
						"0000000000000",--40
						"0000000000000",--41
						"0000000000000",--42
						"0000000000000",--43
						"0000000000000",--44
						"0000000000000",--45
						"0000000000000",--46
						"0000000000000",--47
						"0000000000000",--48
						"0000000000000",--49
						"0001000000001",--50
						"0000010000100",--51
						"0000000000000",--52
						"0000000000000",--53
						"0000000000000",--54
						"0000000000000",--55
						"0000000000000",--56
						"0000000000000",--57
						"0000000000000",--58
						"0000000000000"--59

							
				 );
BEGIN




	

PROCESS(CU_CLK,OPCODE)
VARIABLE X: STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN
IF(STEP="000") THEN  
X:="0000";
ELSE IF(STEP="001") THEN  
X:="0000";
ELSE 
X:=OPCODE;
END IF;
END IF;
ADDRESS<=X&STEP;

IF(CU_CLK'EVENT AND CU_CLK='0') THEN
	CONTROL_BITS<=CONTROL_DATA(CONV_INTEGER(ADDRESS));
	IF(STEP="100") THEN
		STEP<="000";
	ELSE
		STEP<=STEP+1;
	END IF;


	
	

	
END IF;
END PROCESS;
END CONTROL_UNIT;
	
