LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
ENTITY ALU IS 
PORT(
	ALU_CLK: IN STD_LOGIC;
	A: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	B: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	ALU_OUT: IN STD_LOGIC;
	OUTPUT_DATA: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	ARITH_SELECT: IN STD_LOGIC
);
END ALU;

ARCHITECTURE ALU OF ALU IS
BEGIN
PROCESS(ALU_CLK,A,B,ALU_OUT)
VARIABLE ANSWER: SIGNED(7 DOWNTO 0);
VARIABLE OUT_ANSWER: SIGNED(7 DOWNTO 0);
BEGIN
IF(ALU_OUT='1') THEN 
	OUT_ANSWER:=ANSWER;
ELSE IF(ALU_OUT='0') THEN
	OUT_ANSWER:="ZZZZZZZZ";
END IF;
END IF;

IF(ALU_CLK'EVENT AND ALU_CLK='1') THEN
	IF(ARITH_SELECT='1') THEN
	ANSWER:=SIGNED(A)+SIGNED(B);
	ELSE IF (ARITH_SELECT='0') THEN
	ANSWER:=SIGNED(A)- SIGNED(B);
	END IF;

END IF;
OUTPUT_DATA<=STD_LOGIC_VECTOR(OUT_ANSWER);
END IF;

END PROCESS;
END ALU;

	