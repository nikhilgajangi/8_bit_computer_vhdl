	
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY PROGRAM IS
PORT(
	PC_CLK: IN STD_LOGIC;
	PC_OUT: IN STD_LOGIC;
	PC_INC: IN STD_LOGIC;

	PC_ADDRESS: OUT STD_LOGIC_VECTOR( 7 DOWNTO 0)
);
END PROGRAM;


ARCHITECTURE PROGRAM_COUNTER OF PROGRAM IS


BEGIN

PC: PROCESS(PC_CLK,PC_OUT,PC_INC)
VARIABLE PC_BUS: STD_LOGIC_VECTOR(3 DOWNTO 0):="0000";
VARIABLE ADDRESS:STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN
IF(PC_OUT='1') THEN
	ADDRESS:=PC_BUS;
ELSE IF(PC_OUT='0') THEN
	ADDRESS:="ZZZZ";
END IF;
END IF;



IF (PC_CLK'EVENT AND PC_CLK='1') THEN
	IF(PC_INC='1') THEN
		PC_BUS:=PC_BUS+"0001";
	END IF;
PC_ADDRESS<=ADDRESS&"ZZZZ";
END IF;




END PROCESS;
END PROGRAM_COUNTER;